`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: Tristan Richmond
// 
// Create Date: 09/07/2024 12:23:52 PM
// Design Name: 
// Module Name: top_module
// Project Name: 
// Target Devices: Zybo Z7-10
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision: A
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module top_module(

    );
endmodule
